`timescale 1ns / 1ps

module interleaver_tb;

endmodule
